module RRAM();





endmodule
